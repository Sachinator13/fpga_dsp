// cordic.v

// Generated using ACDS version 20.1 720

`timescale 1 ps / 1 ps
module cordic (
		input  wire [15:0] a,      //      a.a
		input  wire        areset, // areset.reset
		output wire [14:0] c,      //      c.c
		input  wire        clk,    //    clk.clk
		output wire [14:0] s       //      s.s
	);

	cordic_CORDIC_0 cordic_0 (
		.clk    (clk),    //    clk.clk
		.areset (areset), // areset.reset
		.a      (a),      //      a.a
		.c      (c),      //      c.c
		.s      (s)       //      s.s
	);

endmodule
